module Condition_Handler(
    input B_instr;
    input [31:26] opcode;
    input flag;  
    input rt; //bits 20:16 de instruction
    output reg  handler_Out;
);


always @* begin


end




endmodule